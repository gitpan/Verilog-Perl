// $Id: v_hier_top2.v 29806 2007-01-10 13:04:28Z wsnyder $
// DESCRIPTION: Verilog-Perl: Example Verilog for testing package
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2000-2007 by Wilson Snyder.

module v_hier_top2 (/*AUTOARG*/
   // Inputs
   clk
   );
   input clk;
endmodule
