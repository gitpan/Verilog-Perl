// $Id: v_hier_noport.v 35110 2007-04-02 13:36:24Z wsnyder $
// DESCRIPTION: Verilog-Perl: Example Verilog for testing package
// This file ONLY is placed into the Public Domain, for any use,
// without warranty, 2000-2007 by Wilson Snyder.

assign foo = 0

module v_hier_noport;
   reg internal;
endmodule
