// $Id: v_hier_top2.v,v 1.2 2001/11/01 21:53:34 wsnyder Exp $
// DESCRIPTION: Verilog-Perl: Example Verilog for testing package

module v_hier_top2 (/*AUTOARG*/
   // Inputs
   clk
   );
   input clk;
endmodule
