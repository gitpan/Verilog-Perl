// $Revision: #3 $$Date: 2002/07/16 $$Author: wsnyder $
// DESCRIPTION: Verilog-Perl: Example Verilog for testing package

module v_hier_top2 (/*AUTOARG*/
   // Inputs
   clk
   );
   input clk;
endmodule
