// $Revision: #1 $$Date: 2002/12/16 $$Author: lab $
// DESCRIPTION: Verilog-Perl: Example Verilog for testing package

module v_hier_top2 (/*AUTOARG*/
   // Inputs
   clk
   );
   input clk;
endmodule
